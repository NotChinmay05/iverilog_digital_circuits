module mux2to1 (
    input  wire sel,
    input  wire [3:0] in0,
    input  wire [3:0] in1,
    output wire [3:0] out
);
    assign out = sel ? in1 : in0;
endmodule
