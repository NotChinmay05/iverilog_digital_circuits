`timescale 1 ns/1 ps
`include "full_adder.v"

module full_adder_tb;

    reg A, B, Cin;
    wire Sum, Cout;

    full_adder uut (.A(A), .B(B), .Cin(Cin), .Sum(Sum), .Cout(Cout));

    initial begin
    $dumpfile("full_adder.vcd");
    $dumpvars(0, full_adder_tb);
        A=0; B=0; Cin=0; #10;
        A=0; B=1; Cin=0; #10;
        A=1; B=0; Cin=0; #10;
        A=1; B=1; Cin=0; #10;

        A=0; B=0; Cin=1; #10;
        A=0; B=1; Cin=1; #10;
        A=1; B=0; Cin=1; #10;
        A=1; B=1; Cin=1; #10;

        #20 $finish;
    end

endmodule
