module jk_ff (
    input J,
    input K,
    input clk,
    output reg Q
);
    initial begin
        Q = 3'b000;
    end
    
    always @(posedge clk) begin
        case ({J, K})
            2'b00: Q <= Q;
            2'b01: Q <= 0;
            2'b10: Q <= 1;
            2'b11: Q <= ~Q;
        endcase
    end

endmodule
